// Definiciones del proyecto MAC
parameter DATA_WIDTH = 16;
parameter ACC_WIDTH  = 40;